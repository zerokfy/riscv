library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        tCYC            : integer := 2
    );
end tb;
